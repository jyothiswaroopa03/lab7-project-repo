//=====================================================================
// Project: 4 core MESI cache design
// File Name: modified_to_invalid_check.sv
// Description: Test for write-miss to D-cache
// Designers: Venky & Suru
//=====================================================================

class modified_to_invalid_check extends base_test;

    //component macro
    `uvm_component_utils(modified_to_invalid_check)

    //Constructor
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction : new

    //UVM build phase
    function void build_phase(uvm_phase phase);
        uvm_config_wrapper::set(this, "tb.vsequencer.run_phase", "default_sequence", modified_to_invalid_check_seq::type_id::get());
        super.build_phase(phase);
    endfunction : build_phase

    //UVM run phase()
    task run_phase(uvm_phase phase);
        `uvm_info(get_type_name(), "Executing modified_to_invalid_check test" , UVM_LOW)
    endtask: run_phase

endclass : modified_to_invalid_check


// Sequence for a Illegal write on I-cache
class modified_to_invalid_check_seq extends base_vseq;
    //object macro
    `uvm_object_utils(modified_to_invalid_check_seq)

    cpu_transaction_c trans;
bit[31:0] addr;
    //constructor
    function new (string name="modified_to_invalid_check_seq");
        super.new(name);
    endfunction : new

    virtual task body();
    repeat(5) begin
`uvm_do_on_with(trans, p_sequencer.cpu_seqr[1], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC;})
addr=trans.address;
        `uvm_do_on_with(trans, p_sequencer.cpu_seqr[0], {request_type == READ_REQ; access_cache_type == DCACHE_ACC; address==addr;})
`uvm_do_on_with(trans, p_sequencer.cpu_seqr[2], {request_type == READ_REQ; access_cache_type == DCACHE_ACC; address==addr;})
`uvm_do_on_with(trans, p_sequencer.cpu_seqr[2], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC; address==addr;})
`uvm_do_on_with(trans, p_sequencer.cpu_seqr[1], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC; address==addr;})


end
    endtask

endclass : modified_to_invalid_check_seq